module schematic1(
	input A,
	input B,
	input C,
	output O10
);


or U5 (O10,A, B, C);

endmodule
