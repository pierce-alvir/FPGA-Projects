module schematic1(
	input A,
	input B,
	output P
);


and U4 (P,A, B);

endmodule
