module schematic1(
	input I3,
	output O4
);


not U2 (O4,I3);

endmodule
